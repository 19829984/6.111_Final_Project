`timescale 1ns / 1ps
`default_nettype none

module trig_lookup #(parameter WIDTH=8) (
    input wire clk_in,
    input wire signed [WIDTH-1:0] angle,
    output logic signed [WIDTH-1:0] cos,
    output logic signed [WIDTH-1:0] sin
);
    always_ff @(posedge clk_in) begin
        case (angle)
			// -1
			8'b11111111: begin
				cos <= 8'b01111111;
				sin <= 8'b11111100;
			end
			// -2
			8'b11111110: begin
				cos <= 8'b01111111;
				sin <= 8'b11111001;
			end
			// -3
			8'b11111101: begin
				cos <= 8'b01111111;
				sin <= 8'b11110110;
			end
			// -4
			8'b11111100: begin
				cos <= 8'b01111111;
				sin <= 8'b11110011;
			end
			// -5
			8'b11111011: begin
				cos <= 8'b01111111;
				sin <= 8'b11110000;
			end
			// -6
			8'b11111010: begin
				cos <= 8'b01111110;
				sin <= 8'b11101101;
			end
			// -7
			8'b11111001: begin
				cos <= 8'b01111110;
				sin <= 8'b11101010;
			end
			// -8
			8'b11111000: begin
				cos <= 8'b01111101;
				sin <= 8'b11100111;
			end
			// -9
			8'b11110111: begin
				cos <= 8'b01111100;
				sin <= 8'b11100011;
			end
			// -10
			8'b11110110: begin
				cos <= 8'b01111100;
				sin <= 8'b11100000;
			end
			// -11
			8'b11110101: begin
				cos <= 8'b01111011;
				sin <= 8'b11011101;
			end
			// -12
			8'b11110100: begin
				cos <= 8'b01111010;
				sin <= 8'b11011010;
			end
			// -13
			8'b11110011: begin
				cos <= 8'b01111001;
				sin <= 8'b11010111;
			end
			// -14
			8'b11110010: begin
				cos <= 8'b01111000;
				sin <= 8'b11010100;
			end
			// -15
			8'b11110001: begin
				cos <= 8'b01110111;
				sin <= 8'b11010001;
			end
			// -16
			8'b11110000: begin
				cos <= 8'b01110110;
				sin <= 8'b11001111;
			end
			// -17
			8'b11101111: begin
				cos <= 8'b01110101;
				sin <= 8'b11001100;
			end
			// -18
			8'b11101110: begin
				cos <= 8'b01110011;
				sin <= 8'b11001001;
			end
			// -19
			8'b11101101: begin
				cos <= 8'b01110010;
				sin <= 8'b11000110;
			end
			// -20
			8'b11101100: begin
				cos <= 8'b01110000;
				sin <= 8'b11000011;
			end
			// -21
			8'b11101011: begin
				cos <= 8'b01101111;
				sin <= 8'b11000000;
			end
			// -22
			8'b11101010: begin
				cos <= 8'b01101101;
				sin <= 8'b10111110;
			end
			// -23
			8'b11101001: begin
				cos <= 8'b01101100;
				sin <= 8'b10111011;
			end
			// -24
			8'b11101000: begin
				cos <= 8'b01101010;
				sin <= 8'b10111000;
			end
			// -25
			8'b11100111: begin
				cos <= 8'b01101000;
				sin <= 8'b10110110;
			end
			// -26
			8'b11100110: begin
				cos <= 8'b01100110;
				sin <= 8'b10110011;
			end
			// -27
			8'b11100101: begin
				cos <= 8'b01100100;
				sin <= 8'b10110001;
			end
			// -28
			8'b11100100: begin
				cos <= 8'b01100010;
				sin <= 8'b10101110;
			end
			// -29
			8'b11100011: begin
				cos <= 8'b01100000;
				sin <= 8'b10101100;
			end
			// -30
			8'b11100010: begin
				cos <= 8'b01011110;
				sin <= 8'b10101010;
			end
			// -31
			8'b11100001: begin
				cos <= 8'b01011100;
				sin <= 8'b10100111;
			end
			// -32
			8'b11100000: begin
				cos <= 8'b01011010;
				sin <= 8'b10100101;
			end
			// -33
			8'b11011111: begin
				cos <= 8'b01011000;
				sin <= 8'b10100011;
			end
			// -34
			8'b11011110: begin
				cos <= 8'b01010101;
				sin <= 8'b10100001;
			end
			// -35
			8'b11011101: begin
				cos <= 8'b01010011;
				sin <= 8'b10011111;
			end
			// -36
			8'b11011100: begin
				cos <= 8'b01010001;
				sin <= 8'b10011101;
			end
			// -37
			8'b11011011: begin
				cos <= 8'b01001110;
				sin <= 8'b10011011;
			end
			// -38
			8'b11011010: begin
				cos <= 8'b01001100;
				sin <= 8'b10011001;
			end
			// -39
			8'b11011001: begin
				cos <= 8'b01001001;
				sin <= 8'b10010111;
			end
			// -40
			8'b11011000: begin
				cos <= 8'b01000111;
				sin <= 8'b10010101;
			end
			// -41
			8'b11010111: begin
				cos <= 8'b01000100;
				sin <= 8'b10010011;
			end
			// -42
			8'b11010110: begin
				cos <= 8'b01000001;
				sin <= 8'b10010010;
			end
			// -43
			8'b11010101: begin
				cos <= 8'b00111111;
				sin <= 8'b10010000;
			end
			// -44
			8'b11010100: begin
				cos <= 8'b00111100;
				sin <= 8'b10001111;
			end
			// -45
			8'b11010011: begin
				cos <= 8'b00111001;
				sin <= 8'b10001101;
			end
			// -46
			8'b11010010: begin
				cos <= 8'b00110110;
				sin <= 8'b10001100;
			end
			// -47
			8'b11010001: begin
				cos <= 8'b00110011;
				sin <= 8'b10001010;
			end
			// -48
			8'b11010000: begin
				cos <= 8'b00110000;
				sin <= 8'b10001001;
			end
			// -49
			8'b11001111: begin
				cos <= 8'b00101110;
				sin <= 8'b10001000;
			end
			// -50
			8'b11001110: begin
				cos <= 8'b00101011;
				sin <= 8'b10000111;
			end
			// -51
			8'b11001101: begin
				cos <= 8'b00101000;
				sin <= 8'b10000110;
			end
			// -52
			8'b11001100: begin
				cos <= 8'b00100101;
				sin <= 8'b10000101;
			end
			// -53
			8'b11001011: begin
				cos <= 8'b00100010;
				sin <= 8'b10000100;
			end
			// -54
			8'b11001010: begin
				cos <= 8'b00011111;
				sin <= 8'b10000011;
			end
			// -55
			8'b11001001: begin
				cos <= 8'b00011100;
				sin <= 8'b10000011;
			end
			// -56
			8'b11001000: begin
				cos <= 8'b00011000;
				sin <= 8'b10000010;
			end
			// -57
			8'b11000111: begin
				cos <= 8'b00010101;
				sin <= 8'b10000001;
			end
			// -58
			8'b11000110: begin
				cos <= 8'b00010010;
				sin <= 8'b10000001;
			end
			// -59
			8'b11000101: begin
				cos <= 8'b00001111;
				sin <= 8'b10000000;
			end
			// -60
			8'b11000100: begin
				cos <= 8'b00001100;
				sin <= 8'b10000000;
			end
			// -61
			8'b11000011: begin
				cos <= 8'b00001001;
				sin <= 8'b10000000;
			end
			// -62
			8'b11000010: begin
				cos <= 8'b00000110;
				sin <= 8'b10000000;
			end
			// -63
			8'b11000001: begin
				cos <= 8'b00000011;
				sin <= 8'b10000000;
			end
			// -64
			8'b11000000: begin
				cos <= 8'b11111111;
				sin <= 8'b10000000;
			end
			// -65
			8'b10111111: begin
				cos <= 8'b11111100;
				sin <= 8'b10000000;
			end
			// -66
			8'b10111110: begin
				cos <= 8'b11111001;
				sin <= 8'b10000000;
			end
			// -67
			8'b10111101: begin
				cos <= 8'b11110110;
				sin <= 8'b10000000;
			end
			// -68
			8'b10111100: begin
				cos <= 8'b11110011;
				sin <= 8'b10000000;
			end
			// -69
			8'b10111011: begin
				cos <= 8'b11110000;
				sin <= 8'b10000000;
			end
			// -70
			8'b10111010: begin
				cos <= 8'b11101101;
				sin <= 8'b10000001;
			end
			// -71
			8'b10111001: begin
				cos <= 8'b11101010;
				sin <= 8'b10000001;
			end
			// -72
			8'b10111000: begin
				cos <= 8'b11100111;
				sin <= 8'b10000010;
			end
			// -73
			8'b10110111: begin
				cos <= 8'b11100011;
				sin <= 8'b10000011;
			end
			// -74
			8'b10110110: begin
				cos <= 8'b11100000;
				sin <= 8'b10000011;
			end
			// -75
			8'b10110101: begin
				cos <= 8'b11011101;
				sin <= 8'b10000100;
			end
			// -76
			8'b10110100: begin
				cos <= 8'b11011010;
				sin <= 8'b10000101;
			end
			// -77
			8'b10110011: begin
				cos <= 8'b11010111;
				sin <= 8'b10000110;
			end
			// -78
			8'b10110010: begin
				cos <= 8'b11010100;
				sin <= 8'b10000111;
			end
			// -79
			8'b10110001: begin
				cos <= 8'b11010001;
				sin <= 8'b10001000;
			end
			// -80
			8'b10110000: begin
				cos <= 8'b11001111;
				sin <= 8'b10001001;
			end
			// -81
			8'b10101111: begin
				cos <= 8'b11001100;
				sin <= 8'b10001010;
			end
			// -82
			8'b10101110: begin
				cos <= 8'b11001001;
				sin <= 8'b10001100;
			end
			// -83
			8'b10101101: begin
				cos <= 8'b11000110;
				sin <= 8'b10001101;
			end
			// -84
			8'b10101100: begin
				cos <= 8'b11000011;
				sin <= 8'b10001111;
			end
			// -85
			8'b10101011: begin
				cos <= 8'b11000000;
				sin <= 8'b10010000;
			end
			// -86
			8'b10101010: begin
				cos <= 8'b10111110;
				sin <= 8'b10010010;
			end
			// -87
			8'b10101001: begin
				cos <= 8'b10111011;
				sin <= 8'b10010011;
			end
			// -88
			8'b10101000: begin
				cos <= 8'b10111000;
				sin <= 8'b10010101;
			end
			// -89
			8'b10100111: begin
				cos <= 8'b10110110;
				sin <= 8'b10010111;
			end
			// -90
			8'b10100110: begin
				cos <= 8'b10110011;
				sin <= 8'b10011001;
			end
			// -91
			8'b10100101: begin
				cos <= 8'b10110001;
				sin <= 8'b10011011;
			end
			// -92
			8'b10100100: begin
				cos <= 8'b10101110;
				sin <= 8'b10011101;
			end
			// -93
			8'b10100011: begin
				cos <= 8'b10101100;
				sin <= 8'b10011111;
			end
			// -94
			8'b10100010: begin
				cos <= 8'b10101010;
				sin <= 8'b10100001;
			end
			// -95
			8'b10100001: begin
				cos <= 8'b10100111;
				sin <= 8'b10100011;
			end
			// -96
			8'b10100000: begin
				cos <= 8'b10100101;
				sin <= 8'b10100101;
			end
			// -97
			8'b10011111: begin
				cos <= 8'b10100011;
				sin <= 8'b10100111;
			end
			// -98
			8'b10011110: begin
				cos <= 8'b10100001;
				sin <= 8'b10101010;
			end
			// -99
			8'b10011101: begin
				cos <= 8'b10011111;
				sin <= 8'b10101100;
			end
			// -100
			8'b10011100: begin
				cos <= 8'b10011101;
				sin <= 8'b10101110;
			end
			// -101
			8'b10011011: begin
				cos <= 8'b10011011;
				sin <= 8'b10110001;
			end
			// -102
			8'b10011010: begin
				cos <= 8'b10011001;
				sin <= 8'b10110011;
			end
			// -103
			8'b10011001: begin
				cos <= 8'b10010111;
				sin <= 8'b10110110;
			end
			// -104
			8'b10011000: begin
				cos <= 8'b10010101;
				sin <= 8'b10111000;
			end
			// -105
			8'b10010111: begin
				cos <= 8'b10010011;
				sin <= 8'b10111011;
			end
			// -106
			8'b10010110: begin
				cos <= 8'b10010010;
				sin <= 8'b10111110;
			end
			// -107
			8'b10010101: begin
				cos <= 8'b10010000;
				sin <= 8'b11000000;
			end
			// -108
			8'b10010100: begin
				cos <= 8'b10001111;
				sin <= 8'b11000011;
			end
			// -109
			8'b10010011: begin
				cos <= 8'b10001101;
				sin <= 8'b11000110;
			end
			// -110
			8'b10010010: begin
				cos <= 8'b10001100;
				sin <= 8'b11001001;
			end
			// -111
			8'b10010001: begin
				cos <= 8'b10001010;
				sin <= 8'b11001100;
			end
			// -112
			8'b10010000: begin
				cos <= 8'b10001001;
				sin <= 8'b11001111;
			end
			// -113
			8'b10001111: begin
				cos <= 8'b10001000;
				sin <= 8'b11010001;
			end
			// -114
			8'b10001110: begin
				cos <= 8'b10000111;
				sin <= 8'b11010100;
			end
			// -115
			8'b10001101: begin
				cos <= 8'b10000110;
				sin <= 8'b11010111;
			end
			// -116
			8'b10001100: begin
				cos <= 8'b10000101;
				sin <= 8'b11011010;
			end
			// -117
			8'b10001011: begin
				cos <= 8'b10000100;
				sin <= 8'b11011101;
			end
			// -118
			8'b10001010: begin
				cos <= 8'b10000011;
				sin <= 8'b11100000;
			end
			// -119
			8'b10001001: begin
				cos <= 8'b10000011;
				sin <= 8'b11100011;
			end
			// -120
			8'b10001000: begin
				cos <= 8'b10000010;
				sin <= 8'b11100111;
			end
			// -121
			8'b10000111: begin
				cos <= 8'b10000001;
				sin <= 8'b11101010;
			end
			// -122
			8'b10000110: begin
				cos <= 8'b10000001;
				sin <= 8'b11101101;
			end
			// -123
			8'b10000101: begin
				cos <= 8'b10000000;
				sin <= 8'b11110000;
			end
			// -124
			8'b10000100: begin
				cos <= 8'b10000000;
				sin <= 8'b11110011;
			end
			// -125
			8'b10000011: begin
				cos <= 8'b10000000;
				sin <= 8'b11110110;
			end
			// -126
			8'b10000010: begin
				cos <= 8'b10000000;
				sin <= 8'b11111001;
			end
			// -127
			8'b10000001: begin
				cos <= 8'b10000000;
				sin <= 8'b11111100;
			end
			// -128
			8'b10000000: begin
				cos <= 8'b10000000;
				sin <= 8'b00000000;
			end
			// 0
			8'b00000000: begin
				cos <= 8'b01111111;
				sin <= 8'b00000000;
			end
			// 1
			8'b00000001: begin
				cos <= 8'b01111111;
				sin <= 8'b00000011;
			end
			// 2
			8'b00000010: begin
				cos <= 8'b01111111;
				sin <= 8'b00000110;
			end
			// 3
			8'b00000011: begin
				cos <= 8'b01111111;
				sin <= 8'b00001001;
			end
			// 4
			8'b00000100: begin
				cos <= 8'b01111111;
				sin <= 8'b00001100;
			end
			// 5
			8'b00000101: begin
				cos <= 8'b01111111;
				sin <= 8'b00001111;
			end
			// 6
			8'b00000110: begin
				cos <= 8'b01111110;
				sin <= 8'b00010010;
			end
			// 7
			8'b00000111: begin
				cos <= 8'b01111110;
				sin <= 8'b00010101;
			end
			// 8
			8'b00001000: begin
				cos <= 8'b01111101;
				sin <= 8'b00011000;
			end
			// 9
			8'b00001001: begin
				cos <= 8'b01111100;
				sin <= 8'b00011100;
			end
			// 10
			8'b00001010: begin
				cos <= 8'b01111100;
				sin <= 8'b00011111;
			end
			// 11
			8'b00001011: begin
				cos <= 8'b01111011;
				sin <= 8'b00100010;
			end
			// 12
			8'b00001100: begin
				cos <= 8'b01111010;
				sin <= 8'b00100101;
			end
			// 13
			8'b00001101: begin
				cos <= 8'b01111001;
				sin <= 8'b00101000;
			end
			// 14
			8'b00001110: begin
				cos <= 8'b01111000;
				sin <= 8'b00101011;
			end
			// 15
			8'b00001111: begin
				cos <= 8'b01110111;
				sin <= 8'b00101110;
			end
			// 16
			8'b00010000: begin
				cos <= 8'b01110110;
				sin <= 8'b00110000;
			end
			// 17
			8'b00010001: begin
				cos <= 8'b01110101;
				sin <= 8'b00110011;
			end
			// 18
			8'b00010010: begin
				cos <= 8'b01110011;
				sin <= 8'b00110110;
			end
			// 19
			8'b00010011: begin
				cos <= 8'b01110010;
				sin <= 8'b00111001;
			end
			// 20
			8'b00010100: begin
				cos <= 8'b01110000;
				sin <= 8'b00111100;
			end
			// 21
			8'b00010101: begin
				cos <= 8'b01101111;
				sin <= 8'b00111111;
			end
			// 22
			8'b00010110: begin
				cos <= 8'b01101101;
				sin <= 8'b01000001;
			end
			// 23
			8'b00010111: begin
				cos <= 8'b01101100;
				sin <= 8'b01000100;
			end
			// 24
			8'b00011000: begin
				cos <= 8'b01101010;
				sin <= 8'b01000111;
			end
			// 25
			8'b00011001: begin
				cos <= 8'b01101000;
				sin <= 8'b01001001;
			end
			// 26
			8'b00011010: begin
				cos <= 8'b01100110;
				sin <= 8'b01001100;
			end
			// 27
			8'b00011011: begin
				cos <= 8'b01100100;
				sin <= 8'b01001110;
			end
			// 28
			8'b00011100: begin
				cos <= 8'b01100010;
				sin <= 8'b01010001;
			end
			// 29
			8'b00011101: begin
				cos <= 8'b01100000;
				sin <= 8'b01010011;
			end
			// 30
			8'b00011110: begin
				cos <= 8'b01011110;
				sin <= 8'b01010101;
			end
			// 31
			8'b00011111: begin
				cos <= 8'b01011100;
				sin <= 8'b01011000;
			end
			// 32
			8'b00100000: begin
				cos <= 8'b01011010;
				sin <= 8'b01011010;
			end
			// 33
			8'b00100001: begin
				cos <= 8'b01011000;
				sin <= 8'b01011100;
			end
			// 34
			8'b00100010: begin
				cos <= 8'b01010101;
				sin <= 8'b01011110;
			end
			// 35
			8'b00100011: begin
				cos <= 8'b01010011;
				sin <= 8'b01100000;
			end
			// 36
			8'b00100100: begin
				cos <= 8'b01010001;
				sin <= 8'b01100010;
			end
			// 37
			8'b00100101: begin
				cos <= 8'b01001110;
				sin <= 8'b01100100;
			end
			// 38
			8'b00100110: begin
				cos <= 8'b01001100;
				sin <= 8'b01100110;
			end
			// 39
			8'b00100111: begin
				cos <= 8'b01001001;
				sin <= 8'b01101000;
			end
			// 40
			8'b00101000: begin
				cos <= 8'b01000111;
				sin <= 8'b01101010;
			end
			// 41
			8'b00101001: begin
				cos <= 8'b01000100;
				sin <= 8'b01101100;
			end
			// 42
			8'b00101010: begin
				cos <= 8'b01000001;
				sin <= 8'b01101101;
			end
			// 43
			8'b00101011: begin
				cos <= 8'b00111111;
				sin <= 8'b01101111;
			end
			// 44
			8'b00101100: begin
				cos <= 8'b00111100;
				sin <= 8'b01110000;
			end
			// 45
			8'b00101101: begin
				cos <= 8'b00111001;
				sin <= 8'b01110010;
			end
			// 46
			8'b00101110: begin
				cos <= 8'b00110110;
				sin <= 8'b01110011;
			end
			// 47
			8'b00101111: begin
				cos <= 8'b00110011;
				sin <= 8'b01110101;
			end
			// 48
			8'b00110000: begin
				cos <= 8'b00110000;
				sin <= 8'b01110110;
			end
			// 49
			8'b00110001: begin
				cos <= 8'b00101110;
				sin <= 8'b01110111;
			end
			// 50
			8'b00110010: begin
				cos <= 8'b00101011;
				sin <= 8'b01111000;
			end
			// 51
			8'b00110011: begin
				cos <= 8'b00101000;
				sin <= 8'b01111001;
			end
			// 52
			8'b00110100: begin
				cos <= 8'b00100101;
				sin <= 8'b01111010;
			end
			// 53
			8'b00110101: begin
				cos <= 8'b00100010;
				sin <= 8'b01111011;
			end
			// 54
			8'b00110110: begin
				cos <= 8'b00011111;
				sin <= 8'b01111100;
			end
			// 55
			8'b00110111: begin
				cos <= 8'b00011100;
				sin <= 8'b01111100;
			end
			// 56
			8'b00111000: begin
				cos <= 8'b00011000;
				sin <= 8'b01111101;
			end
			// 57
			8'b00111001: begin
				cos <= 8'b00010101;
				sin <= 8'b01111110;
			end
			// 58
			8'b00111010: begin
				cos <= 8'b00010010;
				sin <= 8'b01111110;
			end
			// 59
			8'b00111011: begin
				cos <= 8'b00001111;
				sin <= 8'b01111111;
			end
			// 60
			8'b00111100: begin
				cos <= 8'b00001100;
				sin <= 8'b01111111;
			end
			// 61
			8'b00111101: begin
				cos <= 8'b00001001;
				sin <= 8'b01111111;
			end
			// 62
			8'b00111110: begin
				cos <= 8'b00000110;
				sin <= 8'b01111111;
			end
			// 63
			8'b00111111: begin
				cos <= 8'b00000011;
				sin <= 8'b01111111;
			end
			// 64
			8'b01000000: begin
				cos <= 8'b11111111;
				sin <= 8'b01111111;
			end
			// 65
			8'b01000001: begin
				cos <= 8'b11111100;
				sin <= 8'b01111111;
			end
			// 66
			8'b01000010: begin
				cos <= 8'b11111001;
				sin <= 8'b01111111;
			end
			// 67
			8'b01000011: begin
				cos <= 8'b11110110;
				sin <= 8'b01111111;
			end
			// 68
			8'b01000100: begin
				cos <= 8'b11110011;
				sin <= 8'b01111111;
			end
			// 69
			8'b01000101: begin
				cos <= 8'b11110000;
				sin <= 8'b01111111;
			end
			// 70
			8'b01000110: begin
				cos <= 8'b11101101;
				sin <= 8'b01111110;
			end
			// 71
			8'b01000111: begin
				cos <= 8'b11101010;
				sin <= 8'b01111110;
			end
			// 72
			8'b01001000: begin
				cos <= 8'b11100111;
				sin <= 8'b01111101;
			end
			// 73
			8'b01001001: begin
				cos <= 8'b11100011;
				sin <= 8'b01111100;
			end
			// 74
			8'b01001010: begin
				cos <= 8'b11100000;
				sin <= 8'b01111100;
			end
			// 75
			8'b01001011: begin
				cos <= 8'b11011101;
				sin <= 8'b01111011;
			end
			// 76
			8'b01001100: begin
				cos <= 8'b11011010;
				sin <= 8'b01111010;
			end
			// 77
			8'b01001101: begin
				cos <= 8'b11010111;
				sin <= 8'b01111001;
			end
			// 78
			8'b01001110: begin
				cos <= 8'b11010100;
				sin <= 8'b01111000;
			end
			// 79
			8'b01001111: begin
				cos <= 8'b11010001;
				sin <= 8'b01110111;
			end
			// 80
			8'b01010000: begin
				cos <= 8'b11001111;
				sin <= 8'b01110110;
			end
			// 81
			8'b01010001: begin
				cos <= 8'b11001100;
				sin <= 8'b01110101;
			end
			// 82
			8'b01010010: begin
				cos <= 8'b11001001;
				sin <= 8'b01110011;
			end
			// 83
			8'b01010011: begin
				cos <= 8'b11000110;
				sin <= 8'b01110010;
			end
			// 84
			8'b01010100: begin
				cos <= 8'b11000011;
				sin <= 8'b01110000;
			end
			// 85
			8'b01010101: begin
				cos <= 8'b11000000;
				sin <= 8'b01101111;
			end
			// 86
			8'b01010110: begin
				cos <= 8'b10111110;
				sin <= 8'b01101101;
			end
			// 87
			8'b01010111: begin
				cos <= 8'b10111011;
				sin <= 8'b01101100;
			end
			// 88
			8'b01011000: begin
				cos <= 8'b10111000;
				sin <= 8'b01101010;
			end
			// 89
			8'b01011001: begin
				cos <= 8'b10110110;
				sin <= 8'b01101000;
			end
			// 90
			8'b01011010: begin
				cos <= 8'b10110011;
				sin <= 8'b01100110;
			end
			// 91
			8'b01011011: begin
				cos <= 8'b10110001;
				sin <= 8'b01100100;
			end
			// 92
			8'b01011100: begin
				cos <= 8'b10101110;
				sin <= 8'b01100010;
			end
			// 93
			8'b01011101: begin
				cos <= 8'b10101100;
				sin <= 8'b01100000;
			end
			// 94
			8'b01011110: begin
				cos <= 8'b10101010;
				sin <= 8'b01011110;
			end
			// 95
			8'b01011111: begin
				cos <= 8'b10100111;
				sin <= 8'b01011100;
			end
			// 96
			8'b01100000: begin
				cos <= 8'b10100101;
				sin <= 8'b01011010;
			end
			// 97
			8'b01100001: begin
				cos <= 8'b10100011;
				sin <= 8'b01011000;
			end
			// 98
			8'b01100010: begin
				cos <= 8'b10100001;
				sin <= 8'b01010101;
			end
			// 99
			8'b01100011: begin
				cos <= 8'b10011111;
				sin <= 8'b01010011;
			end
			// 100
			8'b01100100: begin
				cos <= 8'b10011101;
				sin <= 8'b01010001;
			end
			// 101
			8'b01100101: begin
				cos <= 8'b10011011;
				sin <= 8'b01001110;
			end
			// 102
			8'b01100110: begin
				cos <= 8'b10011001;
				sin <= 8'b01001100;
			end
			// 103
			8'b01100111: begin
				cos <= 8'b10010111;
				sin <= 8'b01001001;
			end
			// 104
			8'b01101000: begin
				cos <= 8'b10010101;
				sin <= 8'b01000111;
			end
			// 105
			8'b01101001: begin
				cos <= 8'b10010011;
				sin <= 8'b01000100;
			end
			// 106
			8'b01101010: begin
				cos <= 8'b10010010;
				sin <= 8'b01000001;
			end
			// 107
			8'b01101011: begin
				cos <= 8'b10010000;
				sin <= 8'b00111111;
			end
			// 108
			8'b01101100: begin
				cos <= 8'b10001111;
				sin <= 8'b00111100;
			end
			// 109
			8'b01101101: begin
				cos <= 8'b10001101;
				sin <= 8'b00111001;
			end
			// 110
			8'b01101110: begin
				cos <= 8'b10001100;
				sin <= 8'b00110110;
			end
			// 111
			8'b01101111: begin
				cos <= 8'b10001010;
				sin <= 8'b00110011;
			end
			// 112
			8'b01110000: begin
				cos <= 8'b10001001;
				sin <= 8'b00110000;
			end
			// 113
			8'b01110001: begin
				cos <= 8'b10001000;
				sin <= 8'b00101110;
			end
			// 114
			8'b01110010: begin
				cos <= 8'b10000111;
				sin <= 8'b00101011;
			end
			// 115
			8'b01110011: begin
				cos <= 8'b10000110;
				sin <= 8'b00101000;
			end
			// 116
			8'b01110100: begin
				cos <= 8'b10000101;
				sin <= 8'b00100101;
			end
			// 117
			8'b01110101: begin
				cos <= 8'b10000100;
				sin <= 8'b00100010;
			end
			// 118
			8'b01110110: begin
				cos <= 8'b10000011;
				sin <= 8'b00011111;
			end
			// 119
			8'b01110111: begin
				cos <= 8'b10000011;
				sin <= 8'b00011100;
			end
			// 120
			8'b01111000: begin
				cos <= 8'b10000010;
				sin <= 8'b00011000;
			end
			// 121
			8'b01111001: begin
				cos <= 8'b10000001;
				sin <= 8'b00010101;
			end
			// 122
			8'b01111010: begin
				cos <= 8'b10000001;
				sin <= 8'b00010010;
			end
			// 123
			8'b01111011: begin
				cos <= 8'b10000000;
				sin <= 8'b00001111;
			end
			// 124
			8'b01111100: begin
				cos <= 8'b10000000;
				sin <= 8'b00001100;
			end
			// 125
			8'b01111101: begin
				cos <= 8'b10000000;
				sin <= 8'b00001001;
			end
			// 126
			8'b01111110: begin
				cos <= 8'b10000000;
				sin <= 8'b00000110;
			end
			// 127
			8'b01111111: begin
				cos <= 8'b10000000;
				sin <= 8'b00000011;
			end
			// 128
			8'b010000000: begin
				cos <= 8'b10000000;
				sin <= 8'b11111111;
			end
        endcase
    end
endmodule
